// test_sys_top_qsys.v

// Generated using ACDS version 15.0 139

`timescale 1 ps / 1 ps
module test_sys_top_qsys (
		input  wire       clk_50m_clk_in_clk,                      //                   clk_50m_clk_in.clk
		output wire [7:0] led_pio_out8_external_connection_export, // led_pio_out8_external_connection.export
		input  wire       pb_pio_in1_external_connection_export,   //   pb_pio_in1_external_connection.export
		input  wire       reset_0_reset_n,                         //                          reset_0.reset_n
		output wire       temp_lm71cimf_0_conduit_end_cs_n,        //      temp_lm71cimf_0_conduit_end.cs_n
		output wire       temp_lm71cimf_0_conduit_end_sc,          //                                 .sc
		inout  wire       temp_lm71cimf_0_conduit_end_sio          //                                 .sio
	);

	wire  [31:0] master_0_master_readdata;                                  // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                               // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                   // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                      // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                             // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                     // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                 // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [15:0] mm_interconnect_0_temp_lm71cimf_0_avalon_slave_readdata;   // TEMP_LM71CIMF_0:s_readdata -> mm_interconnect_0:TEMP_LM71CIMF_0_avalon_slave_readdata
	wire   [1:0] mm_interconnect_0_temp_lm71cimf_0_avalon_slave_address;    // mm_interconnect_0:TEMP_LM71CIMF_0_avalon_slave_address -> TEMP_LM71CIMF_0:address
	wire         mm_interconnect_0_temp_lm71cimf_0_avalon_slave_read;       // mm_interconnect_0:TEMP_LM71CIMF_0_avalon_slave_read -> TEMP_LM71CIMF_0:s_read
	wire         mm_interconnect_0_temp_lm71cimf_0_avalon_slave_write;      // mm_interconnect_0:TEMP_LM71CIMF_0_avalon_slave_write -> TEMP_LM71CIMF_0:s_write
	wire  [15:0] mm_interconnect_0_temp_lm71cimf_0_avalon_slave_writedata;  // mm_interconnect_0:TEMP_LM71CIMF_0_avalon_slave_writedata -> TEMP_LM71CIMF_0:s_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_0_ocram_1k_s1_chipselect;                  // mm_interconnect_0:ocram_1k_s1_chipselect -> ocram_1k:chipselect
	wire  [31:0] mm_interconnect_0_ocram_1k_s1_readdata;                    // ocram_1k:readdata -> mm_interconnect_0:ocram_1k_s1_readdata
	wire   [7:0] mm_interconnect_0_ocram_1k_s1_address;                     // mm_interconnect_0:ocram_1k_s1_address -> ocram_1k:address
	wire   [3:0] mm_interconnect_0_ocram_1k_s1_byteenable;                  // mm_interconnect_0:ocram_1k_s1_byteenable -> ocram_1k:byteenable
	wire         mm_interconnect_0_ocram_1k_s1_write;                       // mm_interconnect_0:ocram_1k_s1_write -> ocram_1k:write
	wire  [31:0] mm_interconnect_0_ocram_1k_s1_writedata;                   // mm_interconnect_0:ocram_1k_s1_writedata -> ocram_1k:writedata
	wire         mm_interconnect_0_ocram_1k_s1_clken;                       // mm_interconnect_0:ocram_1k_s1_clken -> ocram_1k:clken
	wire         mm_interconnect_0_led_pio_out8_s1_chipselect;              // mm_interconnect_0:led_pio_out8_s1_chipselect -> led_pio_out8:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_out8_s1_readdata;                // led_pio_out8:readdata -> mm_interconnect_0:led_pio_out8_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_out8_s1_address;                 // mm_interconnect_0:led_pio_out8_s1_address -> led_pio_out8:address
	wire         mm_interconnect_0_led_pio_out8_s1_write;                   // mm_interconnect_0:led_pio_out8_s1_write -> led_pio_out8:write_n
	wire  [31:0] mm_interconnect_0_led_pio_out8_s1_writedata;               // mm_interconnect_0:led_pio_out8_s1_writedata -> led_pio_out8:writedata
	wire  [31:0] mm_interconnect_0_pb_pio_in1_s1_readdata;                  // pb_pio_in1:readdata -> mm_interconnect_0:pb_pio_in1_s1_readdata
	wire   [1:0] mm_interconnect_0_pb_pio_in1_s1_address;                   // mm_interconnect_0:pb_pio_in1_s1_address -> pb_pio_in1:address
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [TEMP_LM71CIMF_0:reset, jtag_uart:rst_n, led_pio_out8:reset_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, ocram_1k:reset, pb_pio_in1:reset_n, rst_translator:in_reset, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [ocram_1k:reset_req, rst_translator:reset_req_in]
	wire         master_0_master_reset_reset;                               // master_0:master_reset_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> master_0:clk_reset_reset

	TEMP_LM71CIMF temp_lm71cimf_0 (
		.clk         (clk_50m_clk_in_clk),                                       //   clock_sink.clk
		.reset       (rst_controller_reset_out_reset),                           //   reset_sink.reset
		.address     (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_address),   // avalon_slave.address
		.s_write     (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_write),     //             .write
		.s_writedata (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_writedata), //             .writedata
		.s_read      (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_read),      //             .read
		.s_readdata  (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_readdata),  //             .readdata
		.spi_cs_n    (temp_lm71cimf_0_conduit_end_cs_n),                         //  conduit_end.export
		.spi_sc      (temp_lm71cimf_0_conduit_end_sc),                           //             .export
		.spi_sio     (temp_lm71cimf_0_conduit_end_sio)                           //             .export
	);

	test_sys_top_qsys_jtag_uart jtag_uart (
		.clk            (clk_50m_clk_in_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                                           //               irq.irq
	);

	test_sys_top_qsys_led_pio_out8 led_pio_out8 (
		.clk        (clk_50m_clk_in_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_out8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_out8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_out8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_out8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_out8_s1_readdata),   //                    .readdata
		.out_port   (led_pio_out8_external_connection_export)       // external_connection.export
	);

	test_sys_top_qsys_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_50m_clk_in_clk),                 //          clk.clk
		.clk_reset_reset      (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),            //       master.address
		.master_readdata      (master_0_master_readdata),           //             .readdata
		.master_read          (master_0_master_read),               //             .read
		.master_write         (master_0_master_write),              //             .write
		.master_writedata     (master_0_master_writedata),          //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),        //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),      //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),         //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)         // master_reset.reset
	);

	test_sys_top_qsys_ocram_1k ocram_1k (
		.clk        (clk_50m_clk_in_clk),                       //   clk1.clk
		.address    (mm_interconnect_0_ocram_1k_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ocram_1k_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ocram_1k_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ocram_1k_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ocram_1k_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ocram_1k_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ocram_1k_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)        //       .reset_req
	);

	test_sys_top_qsys_pb_pio_in1 pb_pio_in1 (
		.clk      (clk_50m_clk_in_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pb_pio_in1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pb_pio_in1_s1_readdata), //                    .readdata
		.in_port  (pb_pio_in1_external_connection_export)     // external_connection.export
	);

	test_sys_top_qsys_sysid sysid (
		.clock    (clk_50m_clk_in_clk),                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	test_sys_top_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_50m_clk_clk                                (clk_50m_clk_in_clk),                                        //                              clk_50m_clk.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                            //    jtag_uart_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                        (master_0_master_address),                                   //                          master_0_master.address
		.master_0_master_waitrequest                    (master_0_master_waitrequest),                               //                                         .waitrequest
		.master_0_master_byteenable                     (master_0_master_byteenable),                                //                                         .byteenable
		.master_0_master_read                           (master_0_master_read),                                      //                                         .read
		.master_0_master_readdata                       (master_0_master_readdata),                                  //                                         .readdata
		.master_0_master_readdatavalid                  (master_0_master_readdatavalid),                             //                                         .readdatavalid
		.master_0_master_write                          (master_0_master_write),                                     //                                         .write
		.master_0_master_writedata                      (master_0_master_writedata),                                 //                                         .writedata
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.led_pio_out8_s1_address                        (mm_interconnect_0_led_pio_out8_s1_address),                 //                          led_pio_out8_s1.address
		.led_pio_out8_s1_write                          (mm_interconnect_0_led_pio_out8_s1_write),                   //                                         .write
		.led_pio_out8_s1_readdata                       (mm_interconnect_0_led_pio_out8_s1_readdata),                //                                         .readdata
		.led_pio_out8_s1_writedata                      (mm_interconnect_0_led_pio_out8_s1_writedata),               //                                         .writedata
		.led_pio_out8_s1_chipselect                     (mm_interconnect_0_led_pio_out8_s1_chipselect),              //                                         .chipselect
		.ocram_1k_s1_address                            (mm_interconnect_0_ocram_1k_s1_address),                     //                              ocram_1k_s1.address
		.ocram_1k_s1_write                              (mm_interconnect_0_ocram_1k_s1_write),                       //                                         .write
		.ocram_1k_s1_readdata                           (mm_interconnect_0_ocram_1k_s1_readdata),                    //                                         .readdata
		.ocram_1k_s1_writedata                          (mm_interconnect_0_ocram_1k_s1_writedata),                   //                                         .writedata
		.ocram_1k_s1_byteenable                         (mm_interconnect_0_ocram_1k_s1_byteenable),                  //                                         .byteenable
		.ocram_1k_s1_chipselect                         (mm_interconnect_0_ocram_1k_s1_chipselect),                  //                                         .chipselect
		.ocram_1k_s1_clken                              (mm_interconnect_0_ocram_1k_s1_clken),                       //                                         .clken
		.pb_pio_in1_s1_address                          (mm_interconnect_0_pb_pio_in1_s1_address),                   //                            pb_pio_in1_s1.address
		.pb_pio_in1_s1_readdata                         (mm_interconnect_0_pb_pio_in1_s1_readdata),                  //                                         .readdata
		.sysid_control_slave_address                    (mm_interconnect_0_sysid_control_slave_address),             //                      sysid_control_slave.address
		.sysid_control_slave_readdata                   (mm_interconnect_0_sysid_control_slave_readdata),            //                                         .readdata
		.TEMP_LM71CIMF_0_avalon_slave_address           (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_address),    //             TEMP_LM71CIMF_0_avalon_slave.address
		.TEMP_LM71CIMF_0_avalon_slave_write             (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_write),      //                                         .write
		.TEMP_LM71CIMF_0_avalon_slave_read              (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_read),       //                                         .read
		.TEMP_LM71CIMF_0_avalon_slave_readdata          (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_readdata),   //                                         .readdata
		.TEMP_LM71CIMF_0_avalon_slave_writedata         (mm_interconnect_0_temp_lm71cimf_0_avalon_slave_writedata)   //                                         .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_0_reset_n),                   // reset_in0.reset
		.reset_in1      (master_0_master_reset_reset),        // reset_in1.reset
		.clk            (clk_50m_clk_in_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_0_reset_n),                   // reset_in0.reset
		.reset_in1      (master_0_master_reset_reset),        // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
